`default_nettype none

module MODULENAME(in_wire, out_wire);
    input   wire in_wire;
    output  wire out_wire; 

    assign out_wire = in_wire;
endmodule
